* SKY130 Spice File.
.param
+ sky130_fd_pr__pfet_01v8__lkvth0_diff = .0e-6
+ sky130_fd_pr__pfet_01v8__wlod_diff = .0e-6
+ sky130_fd_pr__pfet_01v8__lku0_diff = 0.0
+ sky130_fd_pr__pfet_01v8__kvsat_diff = 0.5
+ sky130_fd_pr__pfet_01v8__kvth0_diff = 3.29e-8
+ sky130_fd_pr__pfet_01v8__wkvth0_diff = .20e-6
+ sky130_fd_pr__pfet_01v8__ku0_diff = 4.5e-8
+ sky130_fd_pr__pfet_01v8__wku0_diff = .25e-6
