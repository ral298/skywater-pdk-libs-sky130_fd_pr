* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__cap_mim_m3_1 c0 c1 w=1 l=1 mf=1
.param m3_dw = -0.025u
.param tol_m3 = 0.0
.param rm3=0.047
.param rcvia3=3.41
.param tc1rm3= 3.424e-3
.param tc2rm3= -7.739e-7
.param tc1rvia3= 2.366e-3
.param tc2rvia3=-1.025e-5
.param camimc=  2.00e-15
.param cpmimc = 0.19e-15
.param wc = 'w+m3_dw*1e6+tol_m3*1e6'
.param lc = 'l+m3_dw*1e6+tol_m3*1e6'
.param via3_spacing = '(0.17+0.25+0.140)*(0.17+0.25+0.140)'
.param num_contacts = '(wc*lc/via3_spacing)'
.param r1 = 'rm3*(lc)/(wc)'
.param r2 = 'rcvia3/num_contacts'
.param carea = 'camimc*(wc)*(lc)'
.param cperim = 'cpmimc*((wc)+(lc))*2'
.param czero = 'carea + cperim' dev/gauss='0.01*2.8*(carea + cperim)/sqrt(wc*lc*mf)'
c1 c0       a 'czero' tc1 = 0 tc2 = 0.0
rs1 a        b1 'r1' tc1 = {tc1rm3} tc2 = {tc2rm3}
rs2 b1        c1 'r2' tc1 = {tc1rvia3} tc2 = {tc2rvia3}
.ends sky130_fd_pr__cap_mim_m3_1
